library ieee;
use ieee.std_logic_1164.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;


entity top_wrapper is
  port (
    DDR_addr          : inout STD_LOGIC_VECTOR (14 downto 0);
    DDR_ba            : inout STD_LOGIC_VECTOR (2 downto 0);
    DDR_cas_n         : inout STD_LOGIC;
    DDR_ck_n          : inout STD_LOGIC;
    DDR_ck_p          : inout STD_LOGIC;
    DDR_cke           : inout STD_LOGIC;
    DDR_cs_n          : inout STD_LOGIC;
    DDR_dm            : inout STD_LOGIC_VECTOR (3 downto 0);
    DDR_dq            : inout STD_LOGIC_VECTOR (31 downto 0);
    DDR_dqs_n         : inout STD_LOGIC_VECTOR (3 downto 0);
    DDR_dqs_p         : inout STD_LOGIC_VECTOR (3 downto 0);
    DDR_odt           : inout STD_LOGIC;
    DDR_ras_n         : inout STD_LOGIC;
    DDR_reset_n       : inout STD_LOGIC;
    DDR_we_n          : inout STD_LOGIC;
    FIXED_IO_ddr_vrn  : inout STD_LOGIC;
    FIXED_IO_ddr_vrp  : inout STD_LOGIC;
    FIXED_IO_mio      : inout STD_LOGIC_VECTOR (53 downto 0);
    FIXED_IO_ps_clk   : inout STD_LOGIC;
    FIXED_IO_ps_porb  : inout STD_LOGIC;
    FIXED_IO_ps_srstb : inout STD_LOGIC;
    leds              : out   STD_LOGIC_VECTOR(7 downto 0);
    bRight            : in    STD_LOGIC;
    bLeft             : in    STD_LOGIC;
    bDown             : in    STD_LOGIC;
    bUp               : in    STD_LOGIC
  );
end top_wrapper;

architecture STRUCTURE of top_wrapper is
  
  component ps_system is
  port (
    FCLK_CLK0         : out   STD_LOGIC;
    FCLK_RESET0_N     : out   STD_LOGIC;
    DDR_cas_n         : inout STD_LOGIC;
    DDR_cke           : inout STD_LOGIC;
    DDR_ck_n          : inout STD_LOGIC;
    DDR_ck_p          : inout STD_LOGIC;
    DDR_cs_n          : inout STD_LOGIC;
    DDR_reset_n       : inout STD_LOGIC;
    DDR_odt           : inout STD_LOGIC;
    DDR_ras_n         : inout STD_LOGIC;
    DDR_we_n          : inout STD_LOGIC;
    DDR_ba            : inout STD_LOGIC_VECTOR (2 downto 0);
    DDR_addr          : inout STD_LOGIC_VECTOR (14 downto 0);
    DDR_dm            : inout STD_LOGIC_VECTOR (3 downto 0);
    DDR_dq            : inout STD_LOGIC_VECTOR (31 downto 0);
    DDR_dqs_n         : inout STD_LOGIC_VECTOR (3 downto 0);
    DDR_dqs_p         : inout STD_LOGIC_VECTOR (3 downto 0);
    FIXED_IO_mio      : inout STD_LOGIC_VECTOR (53 downto 0);
    FIXED_IO_ddr_vrn  : inout STD_LOGIC;
    FIXED_IO_ddr_vrp  : inout STD_LOGIC;
    FIXED_IO_ps_srstb : inout STD_LOGIC;
    FIXED_IO_ps_clk   : inout STD_LOGIC;
    FIXED_IO_ps_porb  : inout STD_LOGIC;
    bDown             : in    STD_LOGIC;
    bUp               : in    STD_LOGIC
  );
  end component design_1;

  component rModule_leds
    port (
      clk    : in  std_logic;
      rst    : in  std_logic;
      leds   : out std_logic_vector(7 downto 0));
  end component;

  signal FCLK_CLK0     : std_logic;
  signal FCLK_RESET0_N : std_logic;
  signal RESET         : std_logic;
  
begin

  RESET <= not FCLK_RESET0_N;
  
vivado_region : component ps_system
    port map (
      FCLK_CLK0                 => FCLK_CLK0,
      FCLK_RESET0_N             => FCLK_RESET0_N,
      DDR_addr(14 downto 0)     => DDR_addr(14 downto 0),
      DDR_ba(2 downto 0)        => DDR_ba(2 downto 0),
      DDR_cas_n                 => DDR_cas_n,
      DDR_ck_n                  => DDR_ck_n,
      DDR_ck_p                  => DDR_ck_p,
      DDR_cke                   => DDR_cke,
      DDR_cs_n                  => DDR_cs_n,
      DDR_dm(3 downto 0)        => DDR_dm(3 downto 0),
      DDR_dq(31 downto 0)       => DDR_dq(31 downto 0),
      DDR_dqs_n(3 downto 0)     => DDR_dqs_n(3 downto 0),
      DDR_dqs_p(3 downto 0)     => DDR_dqs_p(3 downto 0),
      DDR_odt                   => DDR_odt,
      DDR_ras_n                 => DDR_ras_n,
      DDR_reset_n               => DDR_reset_n,
      DDR_we_n                  => DDR_we_n,
      FIXED_IO_ddr_vrn          => FIXED_IO_ddr_vrn,
      FIXED_IO_ddr_vrp          => FIXED_IO_ddr_vrp,
      FIXED_IO_mio(53 downto 0) => FIXED_IO_mio(53 downto 0),
      FIXED_IO_ps_clk           => FIXED_IO_ps_clk,
      FIXED_IO_ps_porb          => FIXED_IO_ps_porb,
      FIXED_IO_ps_srstb         => FIXED_IO_ps_srstb,
      bDown                     => bDown,
      bUp                       => bUp
    );


rm_leds : rModule_leds
  port map (
    clk    => FCLK_CLK0,
    rst    => RESET,
    leds   => leds);


end STRUCTURE;
