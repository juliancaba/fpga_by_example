`timescale 1 ps / 1 ps

module top_wrapper
(
    leds, 
    DDR_addr,     
    DDR_ba,       
    DDR_cas_n,
    DDR_ck_n,     
    DDR_ck_p,     
    DDR_cke,      
    DDR_cs_n,     
    DDR_dm,       
    DDR_dq,       
    DDR_dqs_n,    
    DDR_dqs_p,    
    DDR_odt,      
    DDR_ras_n,    
    DDR_reset_n,  
    DDR_we_n,     
    FIXED_IO_ddr_vrn,
    FIXED_IO_ddr_vrp, 
    FIXED_IO_mio,
    FIXED_IO_ps_clk,
    FIXED_IO_ps_porb,
    FIXED_IO_ps_srstb
 );
   inout [14:0] DDR_addr;
   inout [2:0] 	DDR_ba;
   inout 	DDR_cas_n;
   inout 	DDR_ck_n;
   inout 	DDR_ck_p;
   inout 	DDR_cke;
   inout 	DDR_cs_n;
   inout [3:0] 	DDR_dm;
   inout [31:0] DDR_dq;
   inout [3:0] 	DDR_dqs_n;
   inout [3:0] 	DDR_dqs_p;
   inout 	DDR_odt;
   inout 	DDR_ras_n;
   inout 	DDR_reset_n;
   inout 	DDR_we_n;
   inout 	FIXED_IO_ddr_vrn;
   inout 	FIXED_IO_ddr_vrp;
   inout [53:0] FIXED_IO_mio;
   inout 	FIXED_IO_ps_clk;
   inout 	FIXED_IO_ps_porb;
   inout 	FIXED_IO_ps_srstb;
   output [7:0] leds;

  wire FCLK_CLK0;
  wire FCLK_RESET0_N;
   
  wire [53:0]FIXED_IO_mio;
  wire FIXED_IO_ps_clk;
  wire FIXED_IO_ps_porb;
  wire FIXED_IO_ps_srstb;
  wire [14:0] DDR_addr;
  wire [2:0] 	DDR_ba;
  wire 	DDR_cas_n;
  wire 	DDR_ck_n;
  wire 	DDR_ck_p;
  wire 	DDR_cke;
  wire 	DDR_cs_n;
  wire [3:0] 	DDR_dm;
  wire [31:0] DDR_dq;
  wire [3:0] 	DDR_dqs_n;
  wire [3:0] 	DDR_dqs_p;
  wire 	DDR_odt;
  wire 	DDR_ras_n;
  wire 	DDR_reset_n;
  wire 	DDR_we_n;
  wire 	FIXED_IO_ddr_vrn;
  wire 	FIXED_IO_ddr_vrp;
   
ps_system vivado_region
       (.FCLK_CLK0(FCLK_CLK0),
	.FCLK_RESET0_N(FCLK_RESET0_N),
	.DDR_cas_n(DDR_cas_n),
	.DDR_cke(DDR_cke),
	.DDR_ck_n(DDR_ck_n),
	.DDR_ck_p(DDR_ck_p),
	.DDR_cs_n(DDR_cs_n),
	.DDR_reset_n(DDR_reset_n),
	.DDR_odt(DDR_odt),
	.DDR_ras_n(DDR_ras_n),
	.DDR_we_n(DDR_we_n),
	.DDR_ba(DDR_ba),
	.DDR_addr(DDR_addr),
	.DDR_dm(DDR_dm),
	.DDR_dq(DDR_dq),
	.DDR_dqs_n(DDR_dqs_n),
	.DDR_dqs_P(DDR_dqs_p),
	.FIXED_IO_ddr_vrn(FIXED_IO_ddr_vrn),
	.FIXED_IO_ddr_vrp(FIXED_IO_ddr_vrp),
        .FIXED_IO_mio(FIXED_IO_mio),
        .FIXED_IO_ps_srstb(FIXED_IO_ps_srstb),	
        .FIXED_IO_ps_clk(FIXED_IO_ps_clk),
        .FIXED_IO_ps_porb(FIXED_IO_ps_porb)
	);

top_reconfig top_dpr
        (.clk(FCLK_CLK0), // 100 MHz clock
         .rst(~FCLK_RESET0_N), // Reset when HIGH
         .leds(leds)); 
        
endmodule // top_wrapper
