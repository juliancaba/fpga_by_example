package readTypes is
  
  type endType is (etNONE, etSIZE, etENDWORD);

end readTypes;
